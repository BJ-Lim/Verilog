module mips_single(clk, reset);
	input clk, reset;
	
	//instruction bus
	wire [31:0] instr;
	
	//break out important fields from instruction
	wire [5:0] opcode, funct;
	wire [4:0] rs, rt, rd, shamt;
	wire [15:0] immed;
	wire [31:0] extend_immed, b_offset;
	wire [25:0] jumpoffset;
	
	assign opcode = instr[31:26];
	assign rs = instr[25:21];
	assign rt = instr[20:16];
	assign rd = instr[15:11];
	assign shamt = instr[10:6];
	assign funct = instr[5:0];
	assign immed = instr[15:0];
	assign jumpoffset = instr[25:0];
	
	//sign-extender
	assign extend_immed = { {16{immed[15]}}, immed };
	
	//branch offset shifter
	assign b_offset = extend_immed << 2;	//address unit is 4bytes.
	
	//datapath signals
	wire [4:0] rfile_wn;
	wire [31:0] rfile_rd1, rfile_rd2, rfile_wd, alu_b, alu_out, b_tgt, pc_next, pc, pc_incr, br_add_out, dmem_rdata;
	
	//control signals
	wire RegWrite, Branch, PCSrc, RegDst, MemtoReg, MemRead, MemWrite, ALUSrc, Zero;
	wire [1:0] ALUOp;
	wire [2:0] Operation;
	
	//module instantiations
	reg32 		PC			(clk, reset, pc_next, pc);
	add32 		PCADD		(pc, 32'd4, pc_incr);
	add32 		BRADD		(pc_incr, b_offset, b_tgt);
	reg_file		RFILE		(clk, RegWrite, rs, rt, rfile_wn, rfile_rd1, rfile_rd2, rfile_wd);
	alu			ALU		(Operation, rfile_rd1, alu_b, alu_out, Zero);
	rom32			IMEM		(pc, instr);
	mem32			DMEM		(clk, MemRead, MemWrite, alu_out, rfile_rd2, dmem_rdata);
	and			BR_AND	(PCSrc, Branch, Zero);
	mux2 #(5)	RFMUX		(RegDst, rt, rd, rfile_wn);
	mux2 #(32)	PCMUX		(PCSrc, pc_incr, b_tgt, pc_next);
	mux2 #(32)	ALUMUX	(ALUSrc, rfile_rd2, extend_immed, alu_b);
	mux2 #(32)	WRMUX		(MemtoReg, alu_out, dmem_rdata, rfile_wd);
	
	
	control_single	CTL	(.opcode(opcode), .RegDst(RegDst), .ALUSrc(ALUSrc), .MemtoReg(MemtoReg),
									.RegWrite(RegWrite), .MemRead(MemRead), .MemWrite(MemWrite), .Branch(Branch),
									.ALUOp(ALUOp));
	alu_ctl		ALUCTL	(ALUOp, funct, Operation);
	
endmodule